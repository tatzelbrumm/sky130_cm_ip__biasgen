** sch_path: /home/cmaier/EDA/efabless/chipalooza2024/sky130_cm_ip__biasgen/xschem/nfet_03v3_gmtest.sch
**.subckt nfet_03v3_gmtest
XM1 Vd Vg GND GND sky130_fd_pr__nfet_03v3_nvt L={l} W={w} nf={nf} ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Evgd Vg Vd Vdref Vd {-egain}
Id net1 Vg {id}
Vdref Vdref GND {vdref}
Vidsense GND net1 0.0
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt



* simulation directives
.option wnflag=1
.option savecurrents
.control
save all
dc Id 10n 10u 10n
plot Vg vs all.Vidsense#branch
*dc vd 0 1.8 0.01 vg 0 1.2 0.1
*plot all.vd1#branch vs D1v8
*plot all.vd2#branch vs D1v8
*save @m.xm1.msky130_fd_pr__nfet_03v3[gm]
*op
write nfet_03v3_gmtest.raw
.endc




.param id     = 10n
.param vdref  = 200m
.param l      = 0.5
.param w      = 1
.param nf     = 1
.param egain  = 1000


**** end user architecture code
**.ends
.GLOBAL GND
.end
