** sch_path: /home/cmaier/EDA/efabless/chipalooza2024/sky130_cm_ip__biasgen/xschem/test_isweep.sch
**.subckt test_isweep
Vdda vdda GND {avdd}
.save i(vdda)
Ibias vdda in {ibias}
Vres res GND {rload}
Bload1 out[1] GND i=(v(out[1])-v(ofs))/v(res)
Vofs ofs GND {vofs}
xDUT vdda vpb vpc out[2] out[1] in GND en[2] en[1] vddd poweron sky130_cm_ip__biasgen l={l} w={w} nf={nf} lc={lc} wc={wc} nfc={nfc}
+ lb={lb} wb={wb} nfb={nfb} ln={lnmos} wn={wnmos} nfn={nfnmos}
Vddd vddd GND {dvdd}
.save i(vddd)
Ven[2] en[2] GND {dvdd}
Ven[1] en[1] GND {dvdd}
.save i(ven[2:1])
* tap: out[2:1] --> out[1]
Bload2 out[2] GND i=(v(out[2])-v(ofs))/v(res)
* tap: out[2:1] --> out[2]
Vpoweron poweron GND {dvdd}
.save i(vpoweron)
**** begin user architecture code

* device parameters
.param l      = 8
.param w      = 2
.param nf     = 1
.param lc     = 0.5
.param wc     = 2
.param nfc    = 1
.param lb     = 18
.param wb     = 1
.param nfb    = 1
.param lnmos  = 8
.param wnmos  = 2
.param nfn    = 1
* instrumentation parameters
.param avdd   = 3.3
.param dvdd   = 1.8
.param ibias  = 50n
.param rload  = 100k
.param vofs   = 1
* simulation parameters
.param celsius = 85
.param imin   = 50n
.param imax   = 1u
.param iinc   = 50n


** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt



* simulation directives
.option wnflag=1
.options gmin=1e-15 abstol=1p
.option savecurrents
.temp {celsius}
.dc Ibias {imin} {imax} {iinc}
.control
save all
run
let Iavg=(@bload1[i]+@bload2[i])/2
let dIio=Iavg-@ibias[current]
let dI=@bload2[i]-@bload1[i]
let dIio_I=dIio/@ibias[current]
let dI_I=dI/Iavg
write test_isweep.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  xschem/sky130_cm_ip__biasgen.sym # of pins=9
** sym_path: /home/cmaier/EDA/efabless/chipalooza2024/sky130_cm_ip__biasgen/xschem/sky130_cm_ip__biasgen.sym
** sch_path: /home/cmaier/EDA/efabless/chipalooza2024/sky130_cm_ip__biasgen/xschem/sky130_cm_ip__biasgen.sch
.subckt sky130_cm_ip__biasgen avdd Vpb Vpc Iout[2] Iout[1] Ibin avss en[2] en[1] dvdd poweron  l=8 w=2 nf=1 lc=0.5 wc=2 nfc=1
+ lb=18 wb=1 nfb=1 lnmos=8 wnmos=2 nfnmos=1
*.iopin avss
*.iopin avdd
*.iopin Ibin
*.iopin Vpb
*.iopin Vpc
*.iopin Iout[2],Iout[1]
*.iopin dvdd
*.iopin en[2],en[1]
*.iopin poweron
xsrc avdd Vpb Vpc Iout[2] Iout[1] Igated avss en[2] en[1] dvdd sky130_cm_sources l={l} w={w} nf={nf} lc={lc} wc={wc} nfc={nfc} lb={lb}
+ wb={wb} nfb={nfb} ln={lnmos} wn={wnmos} nfn={nfnmos}
xpower avdd Vpb Vpc Ibin Igated dvdd poweron avss sky130_cm_poweroff lpt=1 wpt=4 nfpt=1 lnt=1 wnt=2 nfnt=1 lpu=1 wpu=2 nfpu=1
+ lpd=1 wpd=2 nfpd=1
.ends


* expanding   symbol:  xschem/sky130_cm_sources.sym # of pins=8
** sym_path: /home/cmaier/EDA/efabless/chipalooza2024/sky130_cm_ip__biasgen/xschem/sky130_cm_sources.sym
** sch_path: /home/cmaier/EDA/efabless/chipalooza2024/sky130_cm_ip__biasgen/xschem/sky130_cm_sources.sch
.subckt sky130_cm_sources avdd Vpb Vpc Iout[2] Iout[1] Ibin avss en[2] en[1] dvdd  l=8 w=2 nf=1 lc=0.5 wc=2 nfc=1 lb=18 wb=1 nfb=1
+ lnmos=8 wnmos=2 nfnmos=1
*.iopin avss
*.iopin avdd
*.iopin Ibin
*.iopin Vpb
*.iopin Vpc
*.iopin Iout[2],Iout[1]
*.iopin dvdd
*.iopin en[2],en[1]
XMc3 Vpc Vpc avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L={lb} W={wb} nf={nfb} ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMn1 Ibin Ibin avss avss sky130_fd_pr__nfet_g5v0d10v5 L={lnmos} W={wnmos} nf={nfnmos} ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMn2 Vpc Ibin avss avss sky130_fd_pr__nfet_g5v0d10v5 L={lnmos} W={wnmos} nf={nfnmos} ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMn3 Vpb Ibin avss avss sky130_fd_pr__nfet_g5v0d10v5 L={lnmos} W={wnmos} nf={nfnmos} ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
xlvl[2] avdd vgoff[2] dvdd vgon[2] en[2] avss sky130_cm_levelshifter
xlvl[1] avdd vgoff[1] dvdd vgon[1] en[1] avss sky130_cm_levelshifter
x0 avdd avdd Vpb avss Vpc Vpb sky130_cm_sw_psource l={l} w={w} nf={nf} lc={lc} wc={wc} nfc={nfc} lon=.5 won=1 nfon=1 loff=.5 woff=1
+ nfoff=1
xsrc[2] avdd vgoff[2] Vpb vgon[2] Vpc Iout[2] sky130_cm_sw_psource l={l} w={w} nf={nf} lc={lc} wc={wc} nfc={nfc} lon=.5 won=1 nfon=1
+ loff=.5 woff=1 nfoff=1
xsrc[1] avdd vgoff[1] Vpb vgon[1] Vpc Iout[1] sky130_cm_sw_psource l={l} w={w} nf={nf} lc={lc} wc={wc} nfc={nfc} lon=.5 won=1 nfon=1
+ loff=.5 woff=1 nfoff=1
.ends


* expanding   symbol:  xschem/sky130_cm_poweroff.sym # of pins=8
** sym_path: /home/cmaier/EDA/efabless/chipalooza2024/sky130_cm_ip__biasgen/xschem/sky130_cm_poweroff.sym
** sch_path: /home/cmaier/EDA/efabless/chipalooza2024/sky130_cm_ip__biasgen/xschem/sky130_cm_poweroff.sch
.subckt sky130_cm_poweroff avdd Vpb Vpc Ibin Ibout dvdd en avss  lpt=1 wpt=4 nfpt=1 lnt=1 wnt=2 nfnt=1 lpu=1 wpu=2 nfpu=1 lpd=@1
+ wpd=2 nfpd=1
*.iopin avss
*.iopin avdd
*.iopin Ibin
*.iopin Vpb
*.iopin Vpc
*.iopin dvdd
*.iopin en
*.iopin Ibout
XMnpd Ibout off avss avss sky130_fd_pr__nfet_g5v0d10v5 L={lpd} W={wpd} nf={nfpd} ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
xlvl avdd on dvdd off en avss sky130_cm_levelshifter
XMpt Ibout off Ibin avdd sky130_fd_pr__pfet_g5v0d10v5 L={lpt} W={wpt} nf={nfpt} ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMnt Ibout on Ibin avss sky130_fd_pr__nfet_g5v0d10v5 L={lnt} W={wnt} nf={nfnt} ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMpuc Vpc on avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L={lpu} W={wpu} nf={nfpu} ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMpub Vpb on avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L={lpu} W={wpu} nf={nfpu} ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  xschem/sky130_cm_levelshifter.sym # of pins=6
** sym_path: /home/cmaier/EDA/efabless/chipalooza2024/sky130_cm_ip__biasgen/xschem/sky130_cm_levelshifter.sym
** sch_path: /home/cmaier/EDA/efabless/chipalooza2024/sky130_cm_ip__biasgen/xschem/sky130_cm_levelshifter.sch
.subckt sky130_cm_levelshifter avdd Q dvdd Qb A avss
*.iopin avss
*.iopin avdd
*.iopin A
*.iopin dvdd
*.iopin Qb
*.iopin Q
XMnl1 Q ab avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMnl2 Qb abb avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMpl1 Q Qb avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMpl2 Qb Q avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMn1 ab A avss avss sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMp1 ab A dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMn2 abb ab avss avss sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMp2 abb ab dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  xschem/sky130_cm_sw_psource.sym # of pins=6
** sym_path: /home/cmaier/EDA/efabless/chipalooza2024/sky130_cm_ip__biasgen/xschem/sky130_cm_sw_psource.sym
** sch_path: /home/cmaier/EDA/efabless/chipalooza2024/sky130_cm_ip__biasgen/xschem/sky130_cm_sw_psource.sch
.subckt sky130_cm_sw_psource avdd offb Vpb onb Vpc Iout  l=8 w=2 nf=1 lc=0.5 wc=2 nfc=1 lon=.5 won=1 nfon=1 loff=.5 woff=1 nfoff=1
*.iopin avdd
*.iopin Vpb
*.iopin Vpc
*.iopin Iout
*.iopin offb
*.iopin onb
XMc2 Iout vsw vd avdd sky130_fd_pr__pfet_g5v0d10v5 L={lc} W={wc} nf={nfc} ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 vd Vpb avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L={l} W={w} nf={nf} ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMon Vpc onb vsw avdd sky130_fd_pr__pfet_g5v0d10v5 L={lon} W={won} nf={nfon} ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XMoff vsw offb avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L={loff} W={woff} nf={nfoff} ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
