** sch_path: /home/cmaier/EDA/efabless/chipalooza2024/sky130_cm_ip__biasgen/xschem/sky130_cm_ip__biasgen.sch
.subckt sky130_cm_ip__biasgen avdd Vpb Vpc Iout Ibin avss
*.PININFO avss:B avdd:B Ibin:B Vpb:B Vpc:B Iout:B
XMc1 Vpb Vpc vd1 avdd sky130_fd_pr__pfet_g5v0d10v5 L={lc} W={wc} nf={nfc} m=1
XM1 vd1 Vpb avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L={l} W={w} nf={nf} m=1
XMc2 Iout Vpc vd2 avdd sky130_fd_pr__pfet_g5v0d10v5 L={lc} W={wc} nf={nfc} m=1
XM2 vd2 Vpb avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L={l} W={w} nf={nf} m=1
XMc3 Vpc Vpc avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L={lb} W={wb} nf={nfb} m=1
XMn1 Ibin Ibin avss avss sky130_fd_pr__nfet_g5v0d10v5 L={ln} W={wn} nf={nfn} m=1
XMn2 Vpc Ibin avss avss sky130_fd_pr__nfet_g5v0d10v5 L={ln} W={wn} nf={nfn} m=1
XMn3 Vpb Ibin avss avss sky130_fd_pr__nfet_g5v0d10v5 L={ln} W={wn} nf={nfn} m=1
**** begin user architecture code

* device parameters
.param id     = 10n
.param vdref  = 200m
.param l      = 0.15
.param w      = 1
.param nf     = 1
.param lc     = 0.5
.param wc     = 1
.param nfc    = 1
.param lb     = 0.5
.param wb     = 1
.param nfb    = 1
.param ln     = 0.5
.param wn     = 1
.param nfn    = 1
.param egain  = 10000
* simulation parameters
.param imin      = 1n
.param imax      = 10u
.param iinc      = 1n


**** end user architecture code
.ends
.end
