** sch_path: /home/cmaier/EDA/efabless/chipalooza2024/sky130_cm_ip__biasgen/xschem/nfet_01v8_gmtest.sch
**.subckt nfet_01v8_gmtest
Evgd Vg Vd Vdref Vd {-egain}
Id net1 Vg {id}
Vdref Vdref GND {vdref}
Vidsense GND net1 0.0
XM1 Vd Vg GND GND sky130_fd_pr__nfet_01v8 L={l} W=1 nf={nf} ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt



* simulation directives
.option wnflag=1
.option savecurrents
.dc Id {imin} {imax} {iinc} Vdref {vdmin} {vdmax} {vdinc}
.control
save all
run
let gm = deriv(all.Vidsense#branch)/deriv(Vg)
let gm_id = gm/all.Vidsense#branch
plot Vg vs all.Vidsense#branch
plot gm vs all.Vidsense#branch
plot xlog deriv(all.Vidsense#branch)/(deriv(Vg)*all.Vidsense#branch) vs all.Vidsense#branch
write nfet_01v8_gmtest.raw
.endc



* device parameters
.param id     = 10n
.param vdref  = 200m
.param l      = 0.5
.param w      = 1
.param nf     = 1
.param egain  = 1meg
* simulation parameters
.param imin      = 1n
.param imax      = 10u
.param iinc      = 1n
.param vdmin     = 100m
.param vdmax     = 400m
.param vdinc     = 100m


**** end user architecture code
**.ends
.GLOBAL GND
.end
