** sch_path: /home/cmaier/EDA/efabless/chipalooza2024/sky130_cm_ip__biasgen/xschem/sky130_cm_ip__biasgen.sch
.subckt sky130_cm_ip__biasgen vdd vbp vbn vbr vss
*.PININFO vss:B vdd:B vbp:B vbn:B vbr:B
XM10 net3 vbn vres vss sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=4
XM12 vbp vbp vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XM11 vbn vbn vss vss sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM13 net2 vbp vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=4
XM14 net1 vbp vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=2
XM16 vres vbr net5 vss sky130_fd_pr__nfet_01v8 L=20 W=1 nf=1 m=1
XM15 vbr vbr net4 vss sky130_fd_pr__nfet_01v8 L=20 W=1 nf=1 m=1
Vi1 vbp net3 0
.save i(vi1)
Vi4 net2 vbn 0
.save i(vi4)
Viaux net1 vbr 0
.save i(viaux)
XM18 net5 vbr net6 vss sky130_fd_pr__nfet_01v8 L=20 W=1 nf=1 m=1
XM17 net4 vbr net7 vss sky130_fd_pr__nfet_01v8 L=20 W=1 nf=1 m=1
XM20 net6 vbr net9 vss sky130_fd_pr__nfet_01v8 L=20 W=1 nf=1 m=1
XM19 net7 vbr net8 vss sky130_fd_pr__nfet_01v8 L=20 W=1 nf=1 m=1
XM22 net9 vbr vss vss sky130_fd_pr__nfet_01v8 L=20 W=1 nf=1 m=1
XM21 net8 vbr vss vss sky130_fd_pr__nfet_01v8 L=20 W=1 nf=1 m=1
.ends
.end
